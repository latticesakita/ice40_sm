// UART
// 0x00 8'b0000_0000: RO : RBR : Receiver Buffer Register
// 0x00 8'b0000_0000: WO : THR : Transmitter Holding Register
// 0x04 8'b0000_0100: RW : IER : Interrupt Enable Register
// 0x08 8'b0000_1000: RO : IIR : Interrupt Identification register
// 0x0C 8'b0000_1100:      LCR : not supported
// 0x10 8'b0001_0000:      reserved
// 0x14 8'b0001_0100: RO : LSR : Line status register
// 0x18 8'b0001_1000: RO : TXB : Tx fifo available bytes (16bits)
// 0x1C 8'b0001_1100:      reserved
// 0x20 8'b0010_0000: RW : DLR : Divisor LSB (8bits)
// 0x24 8'b0010_0100: RW : DLR : Divisor MSB (8bits)
// 0x28 8'b0010_1000: RW : DLR : Divisor (16bits)
// 0x2C 8'b0010_1100: WO : TMS : Write Timestamp

`define AHBL_IF


module lsc_uart#(
	parameter CLOCK_FREQ = 48000000,
	parameter UART_BAUDRATE = 115200,
	parameter BUFFER_SIZE = "1K" // Tx buffer

)
(
`ifdef AHBL_IF
	input [31:0]	ahbl_haddr_i,	// AHB address
	input [ 2:0]	ahbl_hburst_i,	// unused
	output [31:0]	ahbl_hrdata_o,	// AHB read data
	input [ 2:0]	ahbl_hsize_i,	// unused
	input [ 1:0]	ahbl_htrans_i,	// AHB transfer type
	input [31:0]	ahbl_hwdata_i,	// AHB write data
	input		ahbl_hready_i,	// unused
	output		ahbl_hreadyout_o,	// AHB ready signal
	output		ahbl_hresp_o,	// unused
	input		ahbl_hsel_i,		// AHB select
	input		ahbl_hwrite_i,	// AHB write enable
`else
        input		apb_penable_i, 
        input		apb_psel_i, 
        input		apb_pwrite_i, 
        input	[31:0]	apb_paddr_i, 
        input	[31:0]	apb_pwdata_i, 
        output	[31:0]	apb_prdata_o, 
        output		apb_pslverr_o, 
        output		apb_pready_o,
`endif

	input		i_rxd,
	output reg	o_txd,
	output	reg		int_o,
	input [31:0]    systime_i,

	input		clk,	// data interface, AHBL clock
	input           resetn
);

localparam UART_BAUD_CLK = CLOCK_FREQ/UART_BAUDRATE;

// from timestamp module
reg [7:0] r_hexchar;
reg       r_hexchar_val;

// uart module
reg	[7:0]	i_din;
reg		i_valid;
reg [7:0]	o_dout;
reg      	o_valid;
wire		o_empty;
wire		fifo_full;
wire [15:0]	fifo_available_bytes;
reg [15:0] r_period;
reg		r_rx_int;
reg		r_rx_int_en; // Rx data receive int enable
reg		r_tx_int_en; // Tx fifo empty int enable

// I/F independent signals
reg [31:0]	r_rdata_o;
wire [31:0]     w_wdata_i;
wire [3:0] w_addr;
wire w_re;
wire w_we;
// time stamp related signals
reg [3:0] r_cnt_tms;
wire w_stb_timestamp;
wire w_timestamp_busy;
assign w_timestamp_busy = (w_stb_timestamp||((&r_cnt_tms)==0));

`ifdef AHBL_IF
// AHBL I/F {{{
// AHBL
reg r_we;
reg r_re;
reg [3:0] r_addr;
assign ahbl_hresp_o = 1'b0;
assign w_addr = r_addr; // ahbl_haddr_i[5:2]; // same as LMMI
assign w_re = (ahbl_hsel_i && ahbl_htrans_i[1] && (!ahbl_hwrite_i));
assign w_we = r_we;
assign ahbl_hreadyout_o = ~(r_we|r_re);
assign ahbl_hrdata_o = r_rdata_o;
assign w_wdata_i     = ahbl_hwdata_i;

always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_we <= 0;
		r_re <= 0;
		r_addr <= 0;
	end
	else begin
		r_we <= (ahbl_hsel_i && ahbl_htrans_i[1] &&   ahbl_hwrite_i);
		r_re <= (ahbl_hsel_i && ahbl_htrans_i[1] && (~ahbl_hwrite_i));
		r_addr <= ahbl_haddr_i[5:2];
	end
end

// AHBL I/F }}}
`else
// APB I/F {{{
assign w_addr = apb_paddr_i[5:2];
assign w_re = (apb_psel_i && apb_penable_i && (!apb_pwrite_i));
assign w_we = (apb_psel_i && apb_penable_i && ( apb_pwrite_i));
assign apb_pready_o = 1'b1;
assign apb_prdata_o = r_rdata_o;
assign w_wdata_i = apb_pwdata_i;
// APB I/F }}}
`endif

// I/F independent reg control {{{
// interrupt is only for uart data reception
reg r_valid_d ;
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_valid_d <= 0;
	end
	else begin
		r_valid_d <= o_valid;
	end
end

always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		int_o <= 0;
	end
	else begin
		int_o <= (r_tx_int_en & o_empty) | (r_rx_int_en & r_rx_int);
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_rx_int <= 0;
	end
	else if (!r_rx_int_en) begin
		r_rx_int <= 0;
	end
	else if (w_re) begin
		if(w_addr == 4'h0) begin
			r_rx_int <= 0;
		end
	end
	else begin
		r_rx_int <= r_rx_int | (o_valid & ~r_valid_d);
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_rdata_o <= 32'd0;
	end
	else if (w_re) begin
		if(w_addr == 4'h0) begin // RBR
			r_rdata_o <= {24'd0,o_dout};
		end
		else if(w_addr == 4'h1) begin // IER
			r_rdata_o <= {30'b0,r_tx_int_en,r_rx_int_en};
		end
		else if(w_addr == 4'h2) begin // IIR
			r_rdata_o[31: 8] <= 24'b0;
			r_rdata_o[ 7: 6]  <= 2'b10;
			r_rdata_o[ 5: 3]  <= 3'b000;
			r_rdata_o[ 2: 0]  <= r_rx_int ? 3'b100 : {1'b0,o_empty,1'b0};
		end
		else if(w_addr == 4'h5) begin // LSR 
			r_rdata_o[31: 8] <= 24'b0;
			r_rdata_o[7] <= 1'b0;
			r_rdata_o[6] <= o_empty & (~o_valid);
			r_rdata_o[5] <= o_empty;
			r_rdata_o[4] <= 1'b0; // break condition, not supported
			r_rdata_o[3] <= 1'b0; // framing error, not supported
			r_rdata_o[2] <= 1'b0; // parity error, not supported
			r_rdata_o[1] <= w_timestamp_busy | fifo_full;
			r_rdata_o[0] <= o_valid;
		end
		else if(w_addr == 4'h6) begin // tx fifo available bytes
			r_rdata_o[31:16] <= 16'b0;
			r_rdata_o[15: 0] <=  w_timestamp_busy ? 0 : fifo_available_bytes;
		end
		else if(w_addr == 4'h8) begin
			r_rdata_o[31:8] <= 0;
			r_rdata_o[ 7:0] <= r_period[7:0];
		end
		else if(w_addr == 4'h9) begin
			r_rdata_o[31:8] <= 0;
			r_rdata_o[ 7:0] <= r_period[15:8];
		end
		else if(w_addr == 4'hA) begin
			r_rdata_o[31:16] <= 0;
			r_rdata_o[15:0] <= r_period;
		end
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		i_din <= 0;
		i_valid <= 0;
	end
	else if(w_we && (w_addr == 4'h0)) begin
		i_din <= w_wdata_i[7:0];
		i_valid <= 1;
	end
	else begin
		i_valid <= 0;
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_period <= UART_BAUD_CLK;
	end
	else if(w_we) begin
		if(w_addr == 4'h8) begin
			r_period[7:0] <= w_wdata_i[ 7:0];
		end
		else if(w_addr == 4'h9) begin
			r_period[15:8] <= w_wdata_i[ 7:0];
		end
		else if(w_addr == 4'hA) begin
			r_period[15:0] <= w_wdata_i[15:0];
		end
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_tx_int_en <= 0; // Tx fifo empty int enable
		r_rx_int_en <= 0; // Rx data receive int enable
	end
	else if(w_we) begin
		if(w_addr == 4'h1) begin
			r_tx_int_en <= w_wdata_i[1];
			r_rx_int_en <= w_wdata_i[0];
		end
	end
end
// }}}

// Tx side {{{
localparam TX_FIFO_BITS = 	(BUFFER_SIZE == "4K") ? 12 :
				(BUFFER_SIZE == "2K") ? 11 : 10;
wire		fifo_we;
wire		fifo_rd;
wire	[7:0]	fifo_din;
wire	[7:0]	fifo_dout;
reg		fifo_empty;
reg	[TX_FIFO_BITS -1:0]	fifo_waddr;
reg	[TX_FIFO_BITS -1:0]	fifo_raddr;
reg	[TX_FIFO_BITS -1:0]	fifo_raddr_clk;
reg	[TX_FIFO_BITS -1:0]	fifo_raddr_lat;
reg		r_fifo_empty;
//wire		fifo_full;
wire	[TX_FIFO_BITS -1:0]	fifo_waddr_p1;

reg	[15:0]	tx_period_cnt;
reg	[3:0]	tx_bit_cnt;	// 0: IDLE, 1: Start, 2~9: bit0~7, A:Stop
reg		tx_bit_tick;

always @(posedge clk)
begin
    if(resetn == 1'b0)
	tx_bit_cnt <= 4'b0;
    else if((tx_bit_cnt == 4'b0) && (fifo_empty == 1'b0))
	tx_bit_cnt <= 4'd1;
    else if((tx_bit_cnt == 4'hA) && tx_bit_tick)
	tx_bit_cnt <= 4'd0;
    else if((tx_bit_cnt != 4'b0) && tx_bit_tick)
	tx_bit_cnt <= tx_bit_cnt + 4'd1;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	tx_period_cnt <= 16'b0;
    else if(tx_bit_cnt == 4'b0)
	tx_period_cnt <= 16'b0;
    else if(tx_period_cnt == 16'b0)
	tx_period_cnt <= r_period;
    else
	tx_period_cnt <= tx_period_cnt - 16'd1;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	tx_bit_tick <= 1'b0;
    else if(tx_period_cnt == 16'd1)
	tx_bit_tick <= 1'b1;
    else
	tx_bit_tick <= 1'b0;
end

//assign fifo_rd = ((tx_bit_cnt == 4'hA) && (tx_period_cnt == 16'd1));
assign fifo_rd = ((tx_bit_cnt == 4'h9) && tx_bit_tick);

always @(posedge clk or negedge resetn)
begin
    if(resetn == 1'b0)
	fifo_raddr <= 0;
    else if(fifo_rd)
	fifo_raddr <= fifo_raddr + 1;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	o_txd <= 1'b0;
    else case(tx_bit_cnt)
	4'd1: // start
	    o_txd <= 1'b0;
	4'd2:
	    o_txd <= fifo_dout[0];
	4'd3:
	    o_txd <= fifo_dout[1];
	4'd4:
	    o_txd <= fifo_dout[2];
	4'd5:
	    o_txd <= fifo_dout[3];
	4'd6:
	    o_txd <= fifo_dout[4];
	4'd7:
	    o_txd <= fifo_dout[5];
	4'd8:
	    o_txd <= fifo_dout[6];
	4'd9:
	    o_txd <= fifo_dout[7];
	default: // stop & idle
	    o_txd <= 1'b1;
    endcase
end

always @(posedge clk)
begin
    fifo_raddr_clk <= fifo_raddr;
end

always @(posedge clk or negedge resetn)
begin
    if(resetn == 1'b0)
	fifo_raddr_lat <= 0;
    else if(fifo_raddr_lat != fifo_raddr_clk)
	fifo_raddr_lat <= fifo_raddr_clk;
end

always @(posedge clk or negedge resetn)
begin
    if(resetn == 1'b0)
	r_fifo_empty <= 1'b1;
    else 
	r_fifo_empty <= fifo_raddr_lat == fifo_waddr ;
end

assign fifo_waddr_p1 = fifo_waddr + 1;

assign fifo_we  = ((!fifo_full) && (i_valid | r_hexchar_val));
assign fifo_din = (i_valid) ? i_din : r_hexchar;

always @(posedge clk or negedge resetn)
begin
    if(resetn == 1'b0)
	fifo_waddr <= 0;
    else if(fifo_we)
	fifo_waddr <= fifo_waddr_p1;
end

always @(posedge clk or negedge resetn)
begin
    if(resetn == 1'b0)
	fifo_empty <= 1'b1;
    else
	fifo_empty <= r_fifo_empty;
end

assign o_empty = r_fifo_empty;

assign fifo_full = fifo_raddr_lat == fifo_waddr_p1;
reg [15:0] r_fifo_bytes;
wire [15:0] w_fifo_raddr_16b;
wire [15:0] w_fifo_waddr_16b;
assign w_fifo_raddr_16b[15:TX_FIFO_BITS+1] = 0;
assign w_fifo_raddr_16b[TX_FIFO_BITS] = (fifo_raddr_lat < fifo_waddr_p1);
assign w_fifo_raddr_16b[TX_FIFO_BITS -1:0] = fifo_raddr_lat;
assign w_fifo_waddr_16b[15:TX_FIFO_BITS] = 0;
assign w_fifo_waddr_16b[TX_FIFO_BITS -1:0] = fifo_waddr_p1;
assign fifo_available_bytes = r_fifo_bytes;
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_fifo_bytes <= 0;
	end
	else begin
		r_fifo_bytes <= w_fifo_raddr_16b - w_fifo_waddr_16b ;
	end
end

generate if(BUFFER_SIZE == "4K") 
begin // 4K byte
    dpram4096x8 u_ram4096x8_0 (
	.wr_clk_i   (clk          ),
	.rd_clk_i   (clk      ),
	.wr_clk_en_i(1'b1         ),
	.rd_en_i    (fifo_rd      ),
	.rd_clk_en_i(1'b1         ),
	.wr_en_i    (fifo_we      ),
	.wr_data_i  (fifo_din     ),
	.wr_addr_i  (fifo_waddr   ),
	.rd_addr_i  (fifo_raddr   ),
	.rd_data_o  (fifo_dout    )
    );
end
else if(BUFFER_SIZE == "2K") 
begin // 2K byte
    dpram2048x8 u_ram2048x8_0 (
	.wr_clk_i   (clk          ),
	.rd_clk_i   (clk      ),
	.wr_clk_en_i(1'b1         ),
	.rd_en_i    (fifo_rd      ),
	.rd_clk_en_i(1'b1         ),
	.wr_en_i    (fifo_we      ),
	.wr_data_i  (fifo_din        ),
	.wr_addr_i  (fifo_waddr[10:0]),
	.rd_addr_i  (fifo_raddr[10:0]),
	.rd_data_o  (fifo_dout    )
    );
end
else if(BUFFER_SIZE == "1K") 
begin
    dpram1024x8 u_ram1024x8_0 (
	.wr_clk_i   (clk          ),
	.rd_clk_i   (clk      ),
	.wr_clk_en_i(1'b1         ),
	.rd_en_i    (fifo_rd      ),
	.rd_clk_en_i(1'b1         ),
	.wr_en_i    (fifo_we      ),
	.wr_data_i  (fifo_din        ),
	.wr_addr_i  (fifo_waddr[9:0]),
	.rd_addr_i  (fifo_raddr[9:0]),
	.rd_data_o  (fifo_dout    )
    );
end
else begin // 512 byte
    dpram512x8 u_ram512x8_0 (
	.wr_clk_i   (clk          ),
	.rd_clk_i   (clk      ),
	.wr_clk_en_i(1'b1         ),
	.rd_en_i    (fifo_rd      ),
	.rd_clk_en_i(1'b1         ),
	.wr_en_i    (fifo_we      ),
	.wr_data_i  (fifo_din     ),
	.wr_addr_i  (fifo_waddr[8:0]),
	.rd_addr_i  (fifo_raddr[8:0]),
	.rd_data_o  (fifo_dout    )
    );
end
endgenerate

// Tx side }}}

// Rx side {{{

reg	[15:0]	rx_period_cnt;
reg	[3:0]	rx_bit_cnt;	// 0: IDLE, 1: Start, 2~9: bit0~7, A:Stop
reg		rx_bit_tick;
reg		rx_sample_tick;

reg	[1:0]	rxd_lat;
reg	[7:0]	rxd_shift;

reg		rx_valid_tg;
reg	[1:0]	rx_valid_tg_clk;

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rxd_lat <= 2'b0;
    else 
	rxd_lat <= {rxd_lat[0], i_rxd};
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rxd_shift <= 8'b0;
    else if(rx_sample_tick)
	rxd_shift <= {rxd_lat[0], rxd_shift[7:1]};
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_valid_tg <= 1'b0;
    else if(rx_sample_tick & (rx_bit_cnt == 4'hA))
	rx_valid_tg <= !rx_valid_tg;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	o_dout <= 8'b0;
    else if(rx_sample_tick & (rx_bit_cnt == 4'hA))
	o_dout <= rxd_shift;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_bit_cnt <= 4'b0;
    else if((rx_bit_cnt == 4'b0) && (rxd_lat == 2'b10))
	rx_bit_cnt <= 4'd1;
    else if((rx_bit_cnt == 4'hA) && rx_bit_tick)
	rx_bit_cnt <= 4'd0;
    else if((rx_bit_cnt != 4'b0) && rx_bit_tick)
	rx_bit_cnt <= rx_bit_cnt + 4'd1;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_period_cnt <= 16'b0;
    else if(rx_bit_cnt == 4'b0)
	rx_period_cnt <= 16'b0;
    else if(rx_period_cnt == 16'b0)
	rx_period_cnt <= r_period;
    else
	rx_period_cnt <= rx_period_cnt - 16'd1;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_bit_tick <= 1'b0;
    else if(rx_period_cnt == 16'd1)
	rx_bit_tick <= 1'b1;
    else
	rx_bit_tick <= 1'b0;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_sample_tick <= 1'b0;
    else if(rx_period_cnt == {1'b0, r_period[15:1]})
	rx_sample_tick <= 1'b1;
    else
	rx_sample_tick <= 1'b0;
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	rx_valid_tg_clk <= 2'b0;
    else 
	rx_valid_tg_clk <= {rx_valid_tg_clk[0], rx_valid_tg};
end

always @(posedge clk)
begin
    if(resetn == 1'b0)
	o_valid <= 1'b0;
    else 
	o_valid <= (rx_valid_tg_clk[0] != rx_valid_tg_clk[1]);
end

// Rx side }}}

// Time stamp {{{
function [7:0] HEX2ASCII 
(
   input  [7:0] HEXDATA
);
begin
      case ( HEXDATA )
        8'h80: HEX2ASCII = "0";
        8'h81: HEX2ASCII = "1";
        8'h82: HEX2ASCII = "2";
        8'h83: HEX2ASCII = "3";
        8'h84: HEX2ASCII = "4";
        8'h85: HEX2ASCII = "5";
        8'h86: HEX2ASCII = "6";
        8'h87: HEX2ASCII = "7";
        8'h88: HEX2ASCII = "8";
        8'h89: HEX2ASCII = "9";
        8'h8A: HEX2ASCII = "A";
        8'h8B: HEX2ASCII = "B";
        8'h8C: HEX2ASCII = "C";
        8'h8D: HEX2ASCII = "D";
        8'h8E: HEX2ASCII = "E";
        8'h8F: HEX2ASCII = "F";
	default: HEX2ASCII = HEXDATA;
      endcase
end
endfunction // HEX2ASCII

reg [31:0] r_systime;
reg r_stb_timestamp;
// reg [7:0] r_hexchar;
// reg       r_hexchar_val;
wire [7:0] w_hex;
assign w_stb_timestamp = (w_we && (w_addr ==4'b10_11) && w_wdata_i[0]);
assign w_hex = 
	(r_cnt_tms ==4'b0000) ? {4'b1000,r_systime[31:28]} :
	(r_cnt_tms ==4'b0001) ? {4'b1000,r_systime[27:24]} :
	(r_cnt_tms ==4'b0010) ? {4'b1000,r_systime[23:20]} :
	(r_cnt_tms ==4'b0011) ? {4'b1000,r_systime[19:16]} :
	(r_cnt_tms ==4'b0100) ? {4'b1000,r_systime[15:12]} :
	(r_cnt_tms ==4'b0101) ? {4'b1000,r_systime[11: 8]} :
	(r_cnt_tms ==4'b0110) ? {4'b1000,r_systime[ 7: 4]} :
	(r_cnt_tms ==4'b0111) ? {4'b1000,r_systime[ 3: 0]} :
	(r_cnt_tms ==4'b1000) ? ":" : " ";

always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_systime <= 0;
		r_stb_timestamp <= 0;
	end
	else if(w_stb_timestamp) begin
		r_systime <= systime_i;
		r_stb_timestamp <= 1;
	end
	else begin
		r_stb_timestamp <= 0;
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_cnt_tms <= 4'b1111;
	end
	else if(r_stb_timestamp) begin
		r_cnt_tms <= 4'b0;
	end
	else if(fifo_full) begin
		r_cnt_tms <= r_cnt_tms;
	end
	else if(r_cnt_tms < 4'b1010) begin
		r_cnt_tms <= r_cnt_tms + 1;
	end
	else begin
		r_cnt_tms <= 4'b1111;
	end
end
always @(posedge clk or negedge resetn) begin
	if(!resetn) begin
		r_hexchar     = 8'h00;
		r_hexchar_val = 1'b0;
	end
	else if(r_cnt_tms < 4'b1010) begin
		r_hexchar     = HEX2ASCII(w_hex);
		r_hexchar_val = 1'b1;
	end
	else begin
		r_hexchar     = 8'h00;
		r_hexchar_val = 1'b0;
	end
end

// Time stamp }}}

endmodule

// vim:foldmethod=marker:
//
