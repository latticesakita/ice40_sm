
`timescale 1 ns / 100 ps

module tb;

// GSR GSR_INST (.GSR_N(1'b1));
// PUR PUR_INST (.PUR(1'b1));

parameter FREQ = 12.0;
parameter PERIOD = 1000.0 / FREQ;

reg rstn;
reg clk;

initial begin
	rstn <= 0;
	#100 rstn <= 1;
end
initial begin
	clk = 1'b0;
	forever #(PERIOD/2) clk = ~clk;
end

wire uart_rx;
wire uart_tx;
wire [15:0] led;
wire scl1_io;
wire sda1_io;
wire scl2_io;
wire sda2_io;
wire spi_cs  ;
wire spi_clk ;
wire spi_mosi;
wire spi_miso;

pullup(uart_rx);
pullup(scl1_io);
pullup(sda1_io);
pullup(scl2_io);
pullup(sda2_io);
pullup(led[0]);
pullup(led[1]);
pullup(led[2]);
pullup(led[3]);
pullup(led[4]);
pullup(led[5]);
pullup(led[6]);
pullup(led[7]);
pullup(led[8]);
pullup(led[9]);
pullup(led[10]);
pullup(led[11]);
pullup(led[12]);
pullup(led[13]);
pullup(led[14]);
pullup(led[15]);
pullup(spi_miso);
pullup(spi_mosi);

ice40_sm_top dut (
	//.rstn_i	(rstn),
	//.clk_i	(clk),
	.rxd_i	(uart_rx),
	.txd_o	(uart_tx),
	.led_o	(led[7:0]),
	.scl_io	({scl2_io,scl1_io}),
	.sda_io	({sda2_io,sda1_io}),
	.spi_cs  	(spi_cs  ),
	.spi_clk 	(spi_clk ), 
	.spi_miso	(spi_miso),
	.spi_mosi	(spi_mosi) 
);
// SPI Flash 
spi_flash spi_flash_i (
	.clk		(spi_clk),
	.cs		(spi_cs),
	.miso		(spi_miso),
	.mosi		(spi_mosi)
);
// I2C slave
i2c_slave_tb ov08x (
	.scl(scl1_io),
	.sda(sda1_io),
	.clk(clk)
);



integer code_log;
integer data_log;
integer spram_init_log;

initial begin
	code_log = $fopen("code.log", "w");
	data_log = $fopen("data.log", "w");
	spram_init_log = $fopen("spram_init.log", "w");
end

// ************************
always @(posedge dut.clk_soc or negedge rstn)
	if(dut.spi_sram_we)
		$fwrite(spram_init_log, "%08X\n", dut.spi_sram_din);
 
// ************************
wire [ 1:0] w_instr_htrans     = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HTRANS;
wire [31:0] w_instr_haddr      = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HADDR;
wire [31:0] w_instr_hwdata     = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HWDATA;
wire [31:0] w_instr_hrdata     = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HRDATA;
wire        w_instr_hwrite     = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HWRITE;
wire        w_instr_hready_o   = dut.ice40_sm_inst.cpu_inst_AHBL_M0_INSTR_interconnect_HREADYOUT;
wire        w_instr_ahb_access = w_instr_htrans[1];
reg  [31:0] r_instr_haddr ;
reg  [31:0] r_instr_hwdata;
reg         r_instr_we;
reg         r_instr_re;

always @(posedge dut.clk_soc or negedge rstn) begin
	if(!rstn) begin
		r_instr_we <= 0;
		r_instr_re <= 0;
		r_instr_haddr <= 0;
	end
	else if(w_instr_ahb_access) begin
		r_instr_we <= w_instr_hwrite;
		r_instr_re <= ~w_instr_hwrite;
		r_instr_haddr <= w_instr_haddr;
	end
	else if(w_instr_hready_o) begin
		r_instr_we <= 0;
		r_instr_re <= 0;
	end
end

always @(posedge dut.clk_soc) begin
	if(!w_instr_hready_o) begin
	end
	else if(r_instr_we) begin
		$display(code_log, "%0t: %08X, %08X", $time, 
			r_instr_haddr,
			w_instr_hwdata);
		$fwrite(code_log, "%0t: %08X, %08X, write\n", $time, 
			r_instr_haddr,
			w_instr_hwdata);
	end
	else if(r_instr_re) begin
		$display(code_log, "%0t: %08X, %08X", $time, 
			r_instr_haddr,
			w_instr_hrdata);
		$fwrite(code_log, "%0t: %08X, %08X, read\n", $time, 
			r_instr_haddr,
			w_instr_hrdata);
	end
end
// ************************
wire [ 1:0] w_data_htrans     = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HTRANS;
wire [31:0] w_data_haddr      = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HADDR;
wire [31:0] w_data_hwdata     = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HWDATA;
wire [31:0] w_data_hrdata     = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HRDATA;
wire        w_data_hwrite     = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HWRITE;
wire        w_data_hready_o   = dut.ice40_sm_inst.cpu_inst_AHBL_M1_DATA_interconnect_HREADYOUT;
wire        w_data_ahb_access = w_data_htrans[1];
reg  [31:0] r_data_haddr ;
reg  [31:0] r_data_hwdata;
reg         r_data_we;
reg         r_data_re;

always @(posedge dut.clk_soc or negedge rstn) begin
	if(!rstn) begin
		r_data_we <= 0;
		r_data_re <= 0;
		r_data_haddr <= 0;
	end
	else if(w_data_ahb_access) begin
		r_data_we <= w_data_hwrite;
		r_data_re <= ~w_data_hwrite;
		r_data_haddr <= w_data_haddr;
	end
	else if(w_data_hready_o) begin
		r_data_we <= 0;
		r_data_re <= 0;
	end
end

always @(posedge dut.clk_soc) begin
	if(!w_data_hready_o) begin
	end
	else if(r_data_we) begin
		$display(data_log, "%0t: %08X, %08X", $time, 
			r_data_haddr,
			w_data_hwdata);
		$fwrite(data_log, "%0t: %08X, %08X, write\n", $time, 
			r_data_haddr,
			w_data_hwdata);
	end
	else if(r_data_re) begin
		$display(data_log, "%0t: %08X, %08X", $time, 
			r_data_haddr,
			w_data_hrdata);
		$fwrite(data_log, "%0t: %08X, %08X, read\n", $time, 
			r_data_haddr,
			w_data_hrdata);
	end
end


endmodule
